library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_signed.all;
--use IEEE.std_logic_arith.all;

entity estagio_1 is
	blabla
end estagio_1;

architecture first of estagio_1 is

	blablabla	 

end first;
