-------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : uc_pipeline
-- Author      : Priscilla
-- Company     : x
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\uc_pipeline\uc_pipeline\compile\pipelineTotal.vhd
-- Generated   : Sun Jul  3 12:45:54 2016
-- From        : c:\My_Designs\uc_pipeline\uc_pipeline\src\pipelineTotal.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;


entity pipelineTotal is 
end pipelineTotal;

architecture pipelineTotal of pipelineTotal is

begin

end pipelineTotal;
