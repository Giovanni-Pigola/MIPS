library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_signed.all;
--use IEEE.std_logic_arith.all;

entity estagio_2 is
	port(
	
	
	
	
	
	)
end estagio_2;

architecture estagio2 of estagio_1 is

	blablabla	 

end estagio2;